// Top level module 

module NES (

);

PPU ppu();
CPU cpu();




endmodule 