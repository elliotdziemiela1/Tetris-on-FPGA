module datapath (

);


endmodule 