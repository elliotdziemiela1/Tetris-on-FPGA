// Picture Processing Unit

module PPU (

);





endmodule 